
`ifndef DUMP_LEVEL
`define DUMP_LEVEL 1
`endif

`ifdef DUMP_EN
dump localdump();
`endif